module hello();
    initial begin
        $display("Hello verilator world");
        $finish();
    end
endmodule
